magic
tech sky130A
magscale 1 2
timestamp 1747664904
<< nwell >>
rect -861 -797 861 797
<< mvpmos >>
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
<< mvpdiff >>
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
<< mvpdiffc >>
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
<< mvnsubdiff >>
rect -795 719 795 731
rect -795 685 -687 719
rect 687 685 795 719
rect -795 673 795 685
rect -795 623 -737 673
rect -795 -623 -783 623
rect -749 -623 -737 623
rect 737 623 795 673
rect -795 -673 -737 -623
rect 737 -623 749 623
rect 783 -623 795 623
rect 737 -673 795 -623
rect -795 -685 795 -673
rect -795 -719 -687 -685
rect 687 -719 795 -685
rect -795 -731 795 -719
<< mvnsubdiffcont >>
rect -687 685 687 719
rect -783 -623 -749 623
rect 749 -623 783 623
rect -687 -719 687 -685
<< poly >>
rect -603 581 -503 597
rect -603 547 -587 581
rect -519 547 -503 581
rect -603 500 -503 547
rect -445 581 -345 597
rect -445 547 -429 581
rect -361 547 -345 581
rect -445 500 -345 547
rect -287 581 -187 597
rect -287 547 -271 581
rect -203 547 -187 581
rect -287 500 -187 547
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 500 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 500 129 547
rect 187 581 287 597
rect 187 547 203 581
rect 271 547 287 581
rect 187 500 287 547
rect 345 581 445 597
rect 345 547 361 581
rect 429 547 445 581
rect 345 500 445 547
rect 503 581 603 597
rect 503 547 519 581
rect 587 547 603 581
rect 503 500 603 547
rect -603 -547 -503 -500
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -603 -597 -503 -581
rect -445 -547 -345 -500
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -445 -597 -345 -581
rect -287 -547 -187 -500
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -500
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -500
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -500
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 187 -597 287 -581
rect 345 -547 445 -500
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 345 -597 445 -581
rect 503 -547 603 -500
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 503 -597 603 -581
<< polycont >>
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
<< locali >>
rect -783 685 -687 719
rect 687 685 783 719
rect -783 623 -749 685
rect 749 623 783 685
rect -603 547 -587 581
rect -519 547 -503 581
rect -445 547 -429 581
rect -361 547 -345 581
rect -287 547 -271 581
rect -203 547 -187 581
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect 187 547 203 581
rect 271 547 287 581
rect 345 547 361 581
rect 429 547 445 581
rect 503 547 519 581
rect 587 547 603 581
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 503 -581 519 -547
rect 587 -581 603 -547
rect -783 -685 -749 -623
rect 749 -685 783 -623
rect -783 -719 -687 -685
rect 687 -719 783 -685
<< viali >>
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
<< metal1 >>
rect -599 581 -507 587
rect -599 547 -587 581
rect -519 547 -507 581
rect -599 541 -507 547
rect -441 581 -349 587
rect -441 547 -429 581
rect -361 547 -349 581
rect -441 541 -349 547
rect -283 581 -191 587
rect -283 547 -271 581
rect -203 547 -191 581
rect -283 541 -191 547
rect -125 581 -33 587
rect -125 547 -113 581
rect -45 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 45 581
rect 113 547 125 581
rect 33 541 125 547
rect 191 581 283 587
rect 191 547 203 581
rect 271 547 283 581
rect 191 541 283 547
rect 349 581 441 587
rect 349 547 361 581
rect 429 547 441 581
rect 349 541 441 547
rect 507 581 599 587
rect 507 547 519 581
rect 587 547 599 581
rect 507 541 599 547
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect -599 -547 -507 -541
rect -599 -581 -587 -547
rect -519 -581 -507 -547
rect -599 -587 -507 -581
rect -441 -547 -349 -541
rect -441 -581 -429 -547
rect -361 -581 -349 -547
rect -441 -587 -349 -581
rect -283 -547 -191 -541
rect -283 -581 -271 -547
rect -203 -581 -191 -547
rect -283 -587 -191 -581
rect -125 -547 -33 -541
rect -125 -581 -113 -547
rect -45 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 45 -547
rect 113 -581 125 -547
rect 33 -587 125 -581
rect 191 -547 283 -541
rect 191 -581 203 -547
rect 271 -581 283 -547
rect 191 -587 283 -581
rect 349 -547 441 -541
rect 349 -581 361 -547
rect 429 -581 441 -547
rect 349 -587 441 -581
rect 507 -547 599 -541
rect 507 -581 519 -547
rect 587 -581 599 -547
rect 507 -587 599 -581
<< properties >>
string FIXED_BBOX -766 -702 766 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
