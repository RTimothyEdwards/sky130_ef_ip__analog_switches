magic
tech sky130A
magscale 1 2
timestamp 1747665862
<< metal1 >>
rect 612 -2059 764 -2051
rect 612 -2966 620 -2059
rect 754 -2966 764 -2059
rect 612 -2974 764 -2966
<< via1 >>
rect 620 -2966 754 -2059
<< metal2 >>
rect 612 -2059 764 -2051
rect 612 -2966 620 -2059
rect 754 -2966 764 -2059
rect 612 -2974 764 -2966
<< end >>
