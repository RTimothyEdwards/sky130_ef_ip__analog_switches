magic
tech sky130A
magscale 1 2
timestamp 1747666027
<< pwell >>
rect -673 -414 673 414
<< mvnmos >>
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
<< mvndiff >>
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
<< mvndiffc >>
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
<< mvpsubdiff >>
rect -637 366 637 378
rect -637 332 -529 366
rect 529 332 637 366
rect -637 320 637 332
rect -637 314 -579 320
rect -637 -314 -625 314
rect -591 -314 -579 314
rect 579 314 637 320
rect -637 -320 -579 -314
rect 579 -314 591 314
rect 625 -314 637 314
rect 579 -320 637 -314
rect -637 -332 637 -320
rect -637 -366 -529 -332
rect 529 -366 637 -332
rect -637 -378 637 -366
<< mvpsubdiffcont >>
rect -529 332 529 366
rect -625 -314 -591 314
rect 591 -314 625 314
rect -529 -366 529 -332
<< poly >>
rect -445 272 -345 288
rect -445 238 -429 272
rect -361 238 -345 272
rect -445 200 -345 238
rect -287 272 -187 288
rect -287 238 -271 272
rect -203 238 -187 272
rect -287 200 -187 238
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect 187 272 287 288
rect 187 238 203 272
rect 271 238 287 272
rect 187 200 287 238
rect 345 272 445 288
rect 345 238 361 272
rect 429 238 445 272
rect 345 200 445 238
rect -445 -238 -345 -200
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -445 -288 -345 -272
rect -287 -238 -187 -200
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -287 -288 -187 -272
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
rect 187 -238 287 -200
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 187 -288 287 -272
rect 345 -238 445 -200
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 345 -288 445 -272
<< polycont >>
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
<< locali >>
rect -625 332 -529 366
rect 529 332 625 366
rect -625 314 -591 332
rect 591 314 625 332
rect -445 238 -429 272
rect -361 238 -345 272
rect -287 238 -271 272
rect -203 238 -187 272
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect 187 238 203 272
rect 271 238 287 272
rect 345 238 361 272
rect 429 238 445 272
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 345 -272 361 -238
rect 429 -272 445 -238
rect -625 -332 -591 -314
rect 591 -332 625 -314
rect -625 -366 -529 -332
rect 529 -366 625 -332
<< viali >>
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
<< metal1 >>
rect -441 272 -349 278
rect -441 238 -429 272
rect -361 238 -349 272
rect -441 232 -349 238
rect -283 272 -191 278
rect -283 238 -271 272
rect -203 238 -191 272
rect -283 232 -191 238
rect -125 272 -33 278
rect -125 238 -113 272
rect -45 238 -33 272
rect -125 232 -33 238
rect 33 272 125 278
rect 33 238 45 272
rect 113 238 125 272
rect 33 232 125 238
rect 191 272 283 278
rect 191 238 203 272
rect 271 238 283 272
rect 191 232 283 238
rect 349 272 441 278
rect 349 238 361 272
rect 429 238 441 272
rect 349 232 441 238
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect -441 -238 -349 -232
rect -441 -272 -429 -238
rect -361 -272 -349 -238
rect -441 -278 -349 -272
rect -283 -238 -191 -232
rect -283 -272 -271 -238
rect -203 -272 -191 -238
rect -283 -278 -191 -272
rect -125 -238 -33 -232
rect -125 -272 -113 -238
rect -45 -272 -33 -238
rect -125 -278 -33 -272
rect 33 -238 125 -232
rect 33 -272 45 -238
rect 113 -272 125 -238
rect 33 -278 125 -272
rect 191 -238 283 -232
rect 191 -272 203 -238
rect 271 -272 283 -238
rect 191 -278 283 -272
rect 349 -238 441 -232
rect 349 -272 361 -238
rect 429 -272 441 -238
rect 349 -278 441 -272
<< properties >>
string FIXED_BBOX -608 -393 608 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.5 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
